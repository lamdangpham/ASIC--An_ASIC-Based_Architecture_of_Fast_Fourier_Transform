module mem_input (clk, addr, wr_ena, data) ;
parameter DATA_WIDTH =  32;
input clk;
input wr_ena;
input [11:0] addr;
output [DATA_WIDTH-1:0] data;
reg    [DATA_WIDTH-1:0] data;
always@(posedge clk) begin 
    case(addr)
        0: data <=  32'b0_0000_0000_0000_0000_0000_0000_0000_001;//0
        1: data <=  32'b1_0111_1111_0000_0000_0000_0000_0000_001;//1
        2: data <=  32'b1_0111_1110_0000_0000_0000_0000_0000_010;//0.5
        3: data <=  32'b0_0111_1101_0000_0000_0000_0000_0000_011;//0.25    3e8
        4: data <=  32'b0_0111_1100_0000_0000_0000_0000_0000_100;//0.125   3e0
        5: data <=  32'b0_0111_1011_0000_0000_0000_0000_0000_101;//0.0625   3d8
        6: data <=  32'b0_0000_0000_0000_0000_0000_0000_0000_110;//0
        7: data <=  32'b0_0000_0000_0000_0000_0000_0000_0000_111;//0
        8: data <=  32'b0_0000_0000_0000_0000_0000_0000_0001_000;//0
        default: data <= 0;
    endcase
end

endmodule
